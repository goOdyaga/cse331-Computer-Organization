module heplext(input[15:0] a,output [15:0]b,input c);


or or0(b[0],a[0],c);
or or1(b[1],a[1],c);
or or2(b[2],a[2],c);
or or3(b[3],a[3],c);
or or4(b[4],a[4],c);
or or5(b[5],a[5],c);
or or6(b[6],a[6],c);
or or7(b[7],a[7],c);
or or8(b[8],a[8],c);
or or9(b[9],a[9],c);
or or10(b[10],a[10],c);
or or11(b[11],a[11],c);
or or12(b[12],a[12],c);
or or13(b[13],a[13],c);
or or14(b[14],a[14],c);
or or15(b[15],a[15],c);
endmodule