module muxbitcary(input[31:0] a,input[31:0] b,input select,output [31:0]realres);

wire [31:0]res;
	wire [31:0]resb;
	not not4(selectnot,select);
  
  and and1(res[0], a[0], select);
  and and2(res[1], a[1], select);
  and and3(res[2], a[2], select);
  and and4(res[3], a[3], select);
  and and5(res[4], a[4], select);
  and and6(res[5], a[5], select);
  and and7(res[6], a[6], select);
  and and8(res[7], a[7], select);
  and and9(res[8], a[8], select);
  and and10(res[9], a[9], select);
  and and11(res[10], a[10], select);
  and and12(res[11], a[11], select);
  and and13(res[12], a[12], select);
  and and14(res[13], a[13], select);
  and and15(res[14], a[14], select);
  and and16(res[15], a[15], select);
  and and17(res[16], a[16], select);
  and and18(res[17], a[17], select);
  and and19(res[18], a[18], select);
  and and20(res[19], a[19], select);
  and and21(res[20], a[20], select);
  and and22(res[21], a[21], select);
  and and23(res[22], a[22], select);
  and and24(res[23], a[23], select);
  and and25(res[24], a[24], select);
  and and26(res[25], a[25], select);
  and and27(res[26], a[26], select);
  and and28(res[27], a[27], select);
  and and29(res[28], a[28], select);
  and and30(res[29], a[29], select);
  and and31(res[30], a[30], select);
  and and32(res[31], a[31], select);
  
  and and1b(resb[0], b[0], selectnot);
  and and2b(resb[1], b[1], selectnot);
  and and3b(resb[2], b[2], selectnot);
  and and4b(resb[3], b[3], selectnot);
  and and5b(resb[4], b[4], selectnot);
  and and6b(resb[5], b[5], selectnot);
  and and7b(resb[6], b[6], selectnot);
  and and8b(resb[7], b[7], selectnot);
  and and9b(resb[8], b[8], selectnot);
  and and10b(resb[9], b[9], selectnot);
  and and11b(resb[10], b[10], selectnot);
  and and12b(resb[11], b[11], selectnot);
  and and13b(resb[12], b[12], selectnot);
  and and14b(resb[13], b[13], selectnot);
  and and15b(resb[14], b[14], selectnot);
  and and16b(resb[15], b[15], selectnot);
  and and17b(resb[16], b[16], selectnot);
  and and18b(resb[17], b[17], selectnot);
  and and19b(resb[18], b[18], selectnot);
  and and20b(resb[19], b[19], selectnot);
  and and21b(resb[20], b[20], selectnot);
  and and22b(resb[21], b[21], selectnot);
  and and23b(resb[22], b[22], selectnot);
  and and24b(resb[23], b[23], selectnot);
  and and25b(resb[24], b[24], selectnot);
  and and26b(resb[25], b[25], selectnot);
  and and27b(resb[26], b[26], selectnot);
  and and28b(resb[27], b[27], selectnot);
  and and29b(resb[28], b[28], selectnot);
  and and30b(resb[29], b[29], selectnot);
  and and31b(resb[30], b[30], selectnot);
  and and32b(resb[31], b[31], selectnot);
  
   or or1b(realres[0],    resb[0], res[0]);
  or or2b(realres[1],   resb[1], res[1]);
  or or3b(realres[2],   resb[2], res[2]);
  or or4b(realres[3],   resb[3], res[3]);
  or or5b(realres[4],   resb[4], res[4]);
  or or6b(realres[5],   resb[5], res[5]);
  or or7b(realres[6],   resb[6], res[6]);
  or or8b(realres[7],   resb[7], res[7]);
  or or9b(realres[8],   resb[8], res[8]);
  or or10b(realres[9],  resb[9], res[9] );
  or or11b(realres[10], resb[10], res[10]);
  or or12b(realres[11], resb[11], res[11]);
  or or13b(realres[12], resb[12], res[12]);
  or or14b(realres[13], resb[13], res[13]);
  or or15b(realres[14], resb[14], res[14]);
  or or16b(realres[15], resb[15], res[15]);
  or or17b(realres[16], resb[16], res[16]);
  or or18b(realres[17], resb[17], res[17]);
  or or19b(realres[18], resb[18], res[18]);
  or or20b(realres[19], resb[19], res[19]);
  or or21b(realres[20], resb[20], res[20]);
  or or22b(realres[21], resb[21], res[21]);
  or or23b(realres[22], resb[22], res[22]);
  or or24b(realres[23], resb[23], res[23]);
  or or25b(realres[24], resb[24], res[24]);
  or or26b(realres[25], resb[25], res[25]);
  or or27b(realres[26], resb[26], res[26]);
  or or28b(realres[27], resb[27], res[27]);
  or or29b(realres[28], resb[28], res[28]);
  or or30b(realres[29], resb[29], res[29]);
  or or31b(realres[30], resb[30], res[30]);
  or or32b(realres[31], resb[31], res[31]);


endmodule