module and_with_zero(
  
  output  [31:0] res,input signal
);

  and and1(res[0],1, signal);
  and and2(res[1],1, 0);
  and and3(res[2],1, 0);
  and and4(res[3],1, 0);
  and and5(res[4],1, 0);
  and and6(res[5],1, 0);
  and and7(res[6],1, 0);
  and and8(res[7],1, 0);
  and and9(res[8],1, 0);
  and and10(res[9],1, 0);
  and and11(res[10],1,  0);
  and and12(res[11],1,  0);
  and and13(res[12],1,  0);
  and and14(res[13],1,  0);
  and and15(res[14],1,  0);
  and and16(res[15],1,  0);
  and and17(res[16],1,  0);
  and and18(res[17],1,  0);
  and and19(res[18],1,  0);
  and and20(res[19],1,  0);
  and and21(res[20],1,  0);
  and and22(res[21],1,  0);
  and and23(res[22],1,  0);
  and and24(res[23],1,  0);
  and and25(res[24],1,  0);
  and and26(res[25],1,  0);
  and and27(res[26],1,  0);
  and and28(res[27],1,  0);
  and and29(res[28],1,  0);
  and and30(res[29],1,  0);
  and and31(res[30],1,  0);
  and and32(res[31],1,  0);

endmodule
